c(31)=d(0)+d(1)+d(2)+d(3)+d(4)+d(6)+d(7)+d(8)+d(16)+d(20)+d(22)+d(23)+d(26)+;
c(30)=d(1)+d(2)+d(3)+d(4)+d(5)+d(7)+d(8)+d(9)+d(17)+d(21)+d(23)+d(24)+d(27)+;
c(29)=d(0)+d(2)+d(3)+d(4)+d(5)+d(6)+d(8)+d(9)+d(10)+d(18)+d(22)+d(24)+d(25)+d(28)+;
c(28)=d(1)+d(3)+d(4)+d(5)+d(6)+d(7)+d(9)+d(10)+d(11)+d(19)+d(23)+d(25)+d(26)+d(29)+;
c(27)=d(2)+d(4)+d(5)+d(6)+d(7)+d(8)+d(10)+d(11)+d(12)+d(20)+d(24)+d(26)+d(27)+d(30)+;
c(26)=d(0)+d(3)+d(5)+d(6)+d(7)+d(8)+d(9)+d(11)+d(12)+d(13)+d(21)+d(25)+d(27)+d(28)+d(31)+;
c(25)=d(0)+d(2)+d(3)+d(9)+d(10)+d(12)+d(13)+d(14)+d(16)+d(20)+d(23)+d(28)+d(29)+;
c(24)=d(1)+d(3)+d(4)+d(10)+d(11)+d(13)+d(14)+d(15)+d(17)+d(21)+d(24)+d(29)+d(30)+;
c(23)=d(0)+d(2)+d(4)+d(5)+d(11)+d(12)+d(14)+d(15)+d(16)+d(18)+d(22)+d(25)+d(30)+d(31)+;
c(22)=d(0)+d(2)+d(4)+d(5)+d(7)+d(8)+d(12)+d(13)+d(15)+d(17)+d(19)+d(20)+d(22)+d(31)+;
c(21)=d(0)+d(2)+d(4)+d(5)+d(7)+d(9)+d(13)+d(14)+d(18)+d(21)+d(22)+d(26)+;
c(20)=d(1)+d(3)+d(5)+d(6)+d(8)+d(10)+d(14)+d(15)+d(19)+d(22)+d(23)+d(27)+;
c(19)=d(2)+d(4)+d(6)+d(7)+d(9)+d(11)+d(15)+d(16)+d(20)+d(23)+d(24)+d(28)+;
c(18)=d(0)+d(3)+d(5)+d(7)+d(8)+d(10)+d(12)+d(16)+d(17)+d(21)+d(24)+d(25)+d(29)+;
c(17)=d(0)+d(1)+d(4)+d(6)+d(8)+d(9)+d(11)+d(13)+d(17)+d(18)+d(22)+d(25)+d(26)+d(30)+;
c(16)=d(1)+d(2)+d(5)+d(7)+d(9)+d(10)+d(12)+d(14)+d(18)+d(19)+d(23)+d(26)+d(27)+d(31)+;
c(15)=d(1)+d(4)+d(7)+d(10)+d(11)+d(13)+d(15)+d(16)+d(19)+d(22)+d(23)+d(24)+d(26)+d(27)+d(28)+;
c(14)=d(2)+d(5)+d(8)+d(11)+d(12)+d(14)+d(16)+d(17)+d(20)+d(23)+d(24)+d(25)+d(27)+d(28)+d(29)+;
c(13)=d(0)+d(3)+d(6)+d(9)+d(12)+d(13)+d(15)+d(17)+d(18)+d(21)+d(24)+d(25)+d(26)+d(28)+d(29)+d(30)+;
c(12)=d(0)+d(1)+d(4)+d(7)+d(10)+d(13)+d(14)+d(16)+d(18)+d(19)+d(22)+d(25)+d(26)+d(27)+d(29)+d(30)+d(31)+;
c(11)=d(0)+d(3)+d(4)+d(5)+d(6)+d(7)+d(11)+d(14)+d(15)+d(16)+d(17)+d(19)+d(22)+d(27)+d(28)+d(30)+d(31)+;
c(10)=d(0)+d(2)+d(3)+d(5)+d(12)+d(15)+d(17)+d(18)+d(22)+d(26)+d(28)+d(29)+d(31)+;
c(9)=d(2)+d(7)+d(8)+d(13)+d(18)+d(19)+d(20)+d(22)+d(26)+d(27)+d(29)+d(30)+;
c(8)=d(0)+d(3)+d(8)+d(9)+d(14)+d(19)+d(20)+d(21)+d(23)+d(27)+d(28)+d(30)+d(31)+;
c(7)=d(2)+d(3)+d(6)+d(7)+d(8)+d(9)+d(10)+d(15)+d(16)+d(21)+d(23)+d(24)+d(26)+d(28)+d(29)+d(31)+;
c(6)=d(1)+d(2)+d(6)+d(9)+d(10)+d(11)+d(17)+d(20)+d(23)+d(24)+d(25)+d(26)+d(27)+d(29)+d(30)+;
c(5)=d(2)+d(3)+d(7)+d(10)+d(11)+d(12)+d(18)+d(21)+d(24)+d(25)+d(26)+d(27)+d(28)+d(30)+d(31)+;
c(4)=d(0)+d(1)+d(2)+d(6)+d(7)+d(11)+d(12)+d(13)+d(16)+d(19)+d(20)+d(23)+d(25)+d(27)+d(28)+d(29)+d(31)+;
c(3)=d(0)+d(4)+d(6)+d(12)+d(13)+d(14)+d(16)+d(17)+d(21)+d(22)+d(23)+d(24)+d(28)+d(29)+d(30)+;
c(2)=d(0)+d(1)+d(5)+d(7)+d(13)+d(14)+d(15)+d(17)+d(18)+d(22)+d(23)+d(24)+d(25)+d(29)+d(30)+d(31)+;
c(1)=d(3)+d(4)+d(7)+d(14)+d(15)+d(18)+d(19)+d(20)+d(22)+d(24)+d(25)+d(30)+d(31)+;
c(0)=d(0)+d(1)+d(2)+d(3)+d(5)+d(6)+d(7)+d(15)+d(19)+d(21)+d(22)+d(25)+d(31)+;
